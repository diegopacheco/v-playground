module main

fn main() {
  println('Hello! 1+2=${sum(1,1)} ')
}

fn sum(a int,b int) int {
  return a + b
}