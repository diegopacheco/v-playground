module main

fn test_sum() {
	assert sum(1,2) == 3
}